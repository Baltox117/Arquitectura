module LCDASCII(											//Host Side
	CLK,
	RST_N,
	MP,
																	//LCD Module 16X2
	LCD_ON,														//LCD Power ON/OFF
	LCD_BLON,													//LCD Back Light ON/OFF
	LCD_RW,														//LCD Read/Write Select, 0 = Write, 1 = Read
	LCD_EN,														//LCD Enable
	LCD_RS,														//LCD Command/Data Select, 0 = Command, 1 = Data
	LCD_DATA														//LCD Data bus 8 bits
);																	//Host Side
	input			CLK,RST_N;

////////Agregado///////
	input			[255:0]MP;
///////////////////////

	
//LCD Module 16X2
	output		[7:0]LCD_DATA;								//LCD Data bus 8 bits
	output		LCD_ON;										//LCD Power ON/OFF
	output		LCD_BLON;									//LCD Back Light ON/OFF
	output		LCD_RW;										//LCD Read/Write Select, 0 = Write, 1 = Read
	output		LCD_EN;										//LCD Enable
	output		LCD_RS;										//LCD Command/Data Select, 0 = Command, 1 = Data

//Internal Wires/Registers
	reg			[5:0]LUT_INDEX;
	reg			[8:0]LUT_DATA;
	reg			[7:0]LUT_DATA1;
	reg			[5:0]mLCD_ST;
	reg			[17:0]mDLY;
	reg			mLCD_Start;
	reg			[7:0]mLCD_DATA;
	reg			mLCD_RS;
	wire			mLCD_Done;
	parameter	LCD_INTIAL=0;
	parameter	LCD_LINE1=5;
	parameter	LCD_CH_LINE=LCD_LINE1+16;
	parameter	LCD_LINE2=LCD_LINE1+16+1;
	parameter	LUT_SIZE=LCD_LINE1+32+1;

//LCD ON
	assign		LCD_ON=1'b1;
	assign		LCD_BLON=1'b1;

/////////Comentado/////////	
//	wire			[127:0]MP;
//	assign		MP=128'h0123456789abcdeffedcba9876543210;
/////////Comentado/////////	

	reg			[7:0]CHAR;

	always@(posedge CLK or negedge RST_N)
		begin
			if (!RST_N) begin
				LUT_INDEX<=0;
				mLCD_ST<=0;
				mDLY<=0;
				mLCD_Start<=0;
				mLCD_DATA<=0;
				mLCD_RS<=0;
			end else begin
				if (LUT_INDEX<LUT_SIZE) begin
					case (mLCD_ST)
						0:
							begin
								mLCD_DATA<=LUT_DATA[7:0];
								mLCD_RS<=LUT_DATA[8];
								mLCD_Start<=1;
								mLCD_ST<=1;
							end
						1:
							begin
								if (mLCD_Done) begin
									mLCD_Start<=0;
									mLCD_ST<=2;
								end
							end
						2:
							begin
								if (mDLY<18'h3FFFE)
									mDLY<=mDLY+18'h1;
								else begin
										mDLY<=0;
										mLCD_ST<=3;
								end
							end
						3:
							begin
								LUT_INDEX<=LUT_INDEX+6'h1;
								mLCD_ST<=0;
							end
					endcase
				end
			end
		end

	always														//selecciona el nibble a desplegar del registro
		begin
			case (LUT_INDEX)
//Initial
				LCD_INTIAL+0:LUT_DATA1<=8'h00;
				LCD_INTIAL+1:LUT_DATA1<=8'h00;
				LCD_INTIAL+2:LUT_DATA1<=8'h00;
				LCD_INTIAL+3:LUT_DATA1<=8'h00;
				LCD_INTIAL+4:LUT_DATA1<=8'h00;
//Line 1
				LCD_LINE1+0:LUT_DATA1<={MP[255:248]};       
				LCD_LINE1+1:LUT_DATA1<={MP[247:240]};       
				LCD_LINE1+2:LUT_DATA1<={MP[239:232]};       
				LCD_LINE1+3:LUT_DATA1<={MP[231:224]};       
				LCD_LINE1+4:LUT_DATA1<={MP[223:216]};       
				LCD_LINE1+5:LUT_DATA1<={MP[215:208]};       
				LCD_LINE1+6:LUT_DATA1<={MP[207:200]};       
				LCD_LINE1+7:LUT_DATA1<={MP[199:192]};
				LCD_LINE1+8:LUT_DATA1<={MP[191:184]};
				LCD_LINE1+9:LUT_DATA1<={MP[183:176]};
				LCD_LINE1+10:LUT_DATA1<={MP[175:168]};
				LCD_LINE1+11:LUT_DATA1<={MP[167:160]};
				LCD_LINE1+12:LUT_DATA1<={MP[159:152]};
				LCD_LINE1+13:LUT_DATA1<={MP[151:144]};
				LCD_LINE1+14:LUT_DATA1<={MP[143:136]};
				LCD_LINE1+15:LUT_DATA1<={MP[135:128]};
//Change Line
				LCD_CH_LINE:LUT_DATA1<=8'h00;
//Line 2
				LCD_LINE2+0:LUT_DATA1<={MP[127:120]};
				LCD_LINE2+1:LUT_DATA1<={MP[119:112]};
				LCD_LINE2+2:LUT_DATA1<={MP[111:104]};
				LCD_LINE2+3:LUT_DATA1<={MP[103:96]};
				LCD_LINE2+4:LUT_DATA1<={MP[95:88]};
				LCD_LINE2+5:LUT_DATA1<={MP[87:80]};
				LCD_LINE2+6:LUT_DATA1<={MP[79:72]};
				LCD_LINE2+7:LUT_DATA1<={MP[71:64]};
				LCD_LINE2+8:LUT_DATA1<={MP[63:56]};
				LCD_LINE2+9:LUT_DATA1<={MP[55:48]};
				LCD_LINE2+10:LUT_DATA1<={MP[47:40]};
				LCD_LINE2+11:LUT_DATA1<={MP[39:32]};
				LCD_LINE2+12:LUT_DATA1<={MP[31:24]};
				LCD_LINE2+13:LUT_DATA1<={MP[23:16]};
				LCD_LINE2+14:LUT_DATA1<={MP[15:8]}; 
				LCD_LINE2+15:LUT_DATA1<={MP[7:0]}; 
				default:LUT_DATA1<=8'h00;
			endcase
		end

	always
		begin
//			if(LUT_DATA1<10)
//				CHAR=LUT_DATA1+8'h30;
//			else
//				CHAR=LUT_DATA1+8'h37;
			CHAR = LUT_DATA1;
		end

	always														//Manda a cada posicion del LCD caracter o control
		begin
			case(LUT_INDEX)
//Initial
				LCD_INTIAL+0:LUT_DATA<=9'h038;
				LCD_INTIAL+1:LUT_DATA<=9'h00C;
				LCD_INTIAL+2:LUT_DATA<=9'h001;
				LCD_INTIAL+3:LUT_DATA<=9'h006;
				LCD_INTIAL+4:LUT_DATA<=9'h080;
//Line 1
				LCD_LINE1+0:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+1:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+2:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+3:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+4:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+5:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+6:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+7:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+8:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+9:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+10:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+11:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+12:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+13:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+14:LUT_DATA<={1'b1,CHAR};
				LCD_LINE1+15:LUT_DATA<={1'b1,CHAR};
//Change Line
				LCD_CH_LINE:LUT_DATA<=9'h0C0;
//Line 2
				LCD_LINE2+0:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+1:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+2:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+3:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+4:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+5:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+6:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+7:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+8:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+9:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+10:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+11:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+12:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+13:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+14:LUT_DATA<={1'b1,CHAR};
				LCD_LINE2+15:LUT_DATA<={1'b1,CHAR};
				default:LUT_DATA<=9'h000;
			endcase
		end
		LCD_ControllerASCII u0(									//Host Side
			.iDATA(mLCD_DATA),
			.iRS(mLCD_RS),
			.iStart(mLCD_Start),
			.oDone(mLCD_Done),
			.CLK(CLK),
			.RST_N(RST_N),
//LCD Interface
			.LCD_DATA(LCD_DATA),
			.LCD_RW(LCD_RW),
			.LCD_EN(LCD_EN),
			.LCD_RS(LCD_RS)
		);
endmodule

module LCD_ControllerASCII(										//Host Side
	iDATA,iRS,
	iStart,oDone,
	CLK,RST_N,
//	LCD Interface
	LCD_DATA,
	LCD_RW,
	LCD_EN,
	LCD_RS
);
//CLK
	parameter	CLK_Divide=16;
//Host Side
	input			[7:0]iDATA;
	input			iRS,iStart;
	input			CLK,RST_N;
	output reg	oDone;
//LCD Interface
	output		[7:0]LCD_DATA;
	output reg	LCD_EN;
	output		LCD_RW;
	output		LCD_RS;
//Internal Register
	reg			[4:0]Cont;
	reg			[1:0]ST;
	reg			preStart,mStart;
/////////////////////////////////////////////
//Only write to LCD, bypass iRS to LCD_RS
	assign		LCD_DATA=iDATA; 
	assign		LCD_RW=1'b0;
	assign		LCD_RS=iRS;
/////////////////////////////////////////////
	always@(posedge CLK or negedge RST_N)
		begin
			if (!RST_N) begin
				oDone<=1'b0;
				LCD_EN<=1'b0;
				preStart<=1'b0;
				mStart<=1'b0;
				Cont<=0;
				ST<=0;
			end else	begin
//////Input Start Detect ///////
				preStart<=iStart;
				if ({preStart,iStart}==2'b01) begin
					mStart<=1'b1;
					oDone<=1'b0;
				end
//////////////////////////////////
				if (mStart) begin
					case(ST)
						0:	ST<=1;								//Wait Setup
						1:
							begin
								LCD_EN<=1'b1;
								ST<=2;
							end
						2:
							begin
								if (Cont<CLK_Divide)
									Cont<=Cont+5'h1;
								else
									ST<=3;
							end
						3:
							begin
								LCD_EN<=1'b0;
								mStart<=1'b0;
								oDone<=1'b1;
								Cont<=0;
								ST<=0;
							end
					endcase
				end
			end
		end
endmodule 